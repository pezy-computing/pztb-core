`ifndef PZVIP_TILELINK_DEFINES_SVH
`define PZVIP_TILELINK_DEFINES_SVH

`ifndef PZVIP_TILELINK_MAX_DATA_WIDTH
  `define PZVIP_TILELINK_MAX_DATA_WIDTH 256
`endif

`ifndef PZVIP_TILELINK_MAX_ADDRESS_WIDTH
  `define PZVIP_TILELINK_MAX_ADDRESS_WIDTH  48
`endif

`ifndef PZVIP_TILELINK_MAX_SIZE
  `define PZVIP_TILELINK_MAX_SIZE (2**15)
`endif

`ifndef PZVIP_TILELINK_MAX_ID_WIDTH
  `define PZVIP_TILELINK_MAX_ID_WIDTH 8
`endif

`endif
