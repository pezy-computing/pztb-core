class pzvip_i2c_status extends tue_status;
  `tue_object_default_constructor(pzvip_i2c_status)
  `uvm_object_utils(pzvip_i2c_status)
endclass
