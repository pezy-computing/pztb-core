class pzvip_uart_configuration extends tue_configuration;
  pzvip_uart_vif    vif;
  `tue_object_default_constructor(pzvip_uart_configuration)
  `uvm_object_utils(pzvip_uart_configuration)
endclass
