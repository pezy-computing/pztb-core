class pzvip_spi_status extends tue_status;
  `tue_object_default_constructor(pzvip_spi_status)
  `uvm_object_utils(pzvip_spi_status)
endclass
