`ifndef PZVIP_STREAM_DEFINES_SVH
`define PZVIP_STREAM_DEFINES_SVH

`ifndef PZVIP_STREAM_MAX_DATA_WIDTH
  `define PZVIP_STREAM_MAX_DATA_WIDTH 256
`endif

`endif
