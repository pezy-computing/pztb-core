`ifndef PZVIP_COREBUS_INTERNAL_MACROS_SVH
`define PZVIP_COREBUS_INTERNAL_MACROS_SVH

`define pzvip_corebus_get_mask(WIDTH) ((1 << WIDTH) - 1)

`endif
