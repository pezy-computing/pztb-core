package pzvip_corebus_sample_pkg;
  import  uvm_pkg::*;
  import  tue_pkg::*;
  import  pzvip_corebus_types_pkg::*;
  import  pzvip_corebus_pkg::*;

  `include  "uvm_macros.svh"
  `include  "tue_macros.svh"

  `include  "pzvip_corebus_sample_configuration.svh"
  `include  "pzvip_corebus_sample_write_read_sequence.svh"
  `include  "pzvip_corebus_sample_test.svh"
endpackage
