typedef tue_status_dummy  pzvip_stream_status;
