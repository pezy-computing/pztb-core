class pzvip_uart_status extends tue_status;
  `tue_object_default_constructor(pzvip_uart_status)
  `uvm_object_utils(pzvip_uart_status)
endclass
