//========================================
//
// Copyright (c) 2023 PEZY Computing, K.K.
//                    All Rights Reserved.
//
//========================================
package pztb_pkg;
  typedef enum logic [1:0] {
    PZTB_MEM_INIT_X,
    PZTB_MEM_INIT_0,
    PZTB_MEM_INIT_1,
    PZTB_MEM_INIT_RANDOM
  } pztb_mem_init;
endpackage
